module tempMemory #(
    parameter int SIZE = 8192,
    parameter int N = 13  // log2(SIZE)
)(
    input  logic         clk,
    input  logic         rst,
    input  logic         write_en,
    input  logic [N-1:0] addr,
    input  logic [7:0]   data_in,
    output logic [7:0]   data_out
);

    logic [7:0] mem_array [0:SIZE-1];

    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            int i;
            for (i = 0; i < SIZE; i++) begin
                mem_array[i] <= 8'd0;
            end
        end
        else if (write_en) begin
            mem_array[addr] <= data_in;
        end
    end

    assign data_out = mem_array[addr];

endmodule
